typedef struct packed {
    logic [23:0] I;
    logic [23:0] Q;
} Samp;

typedef struct packed {
    logic [26:0] I;
    logic [26:0] Q;
} Coef;